///////////////////////////////////////////////////////////////////////////////
// Author: Will Chen
//
// Description:
//    * Source file include list for computer vision edge detector testbench
///////////////////////////////////////////////////////////////////////////////


// Testbench source files
`include "verif/tb.sv"  // Manual testbench

