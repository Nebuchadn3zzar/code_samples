initial begin
   $dumpfile("waves.vcd");
   $dumpvars();
   $dumpon();
end

